module datapath(input logic[15:0] X,
                output logic [15:0] answer);

endmodule // datapath
